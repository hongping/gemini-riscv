module helloworld();
    initial begin
        $display("hello");
    end
endmodule